library verilog;
use verilog.vl_types.all;
entity MaquinaSalgados_vlg_vec_tst is
end MaquinaSalgados_vlg_vec_tst;
